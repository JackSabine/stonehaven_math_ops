`include "multiplier_basic_test.sv"
